// TimerSoC.v

// Generated using ACDS version 18.1 625

`timescale 1 ps / 1 ps
module TimerSoC (
		input  wire [1:0]  buttons_export,  //  buttons.export
		input  wire        clk_clk,         //      clk.clk
		output wire [31:0] displays_export, // displays.export
		input  wire [7:0]  gpio_in_export,  //  gpio_in.export
		output wire [7:0]  gpio_out_export, // gpio_out.export
		output wire [9:0]  leds_export,     //     leds.export
		input  wire        reset_reset_n,   //    reset.reset_n
		input  wire [1:0]  switches_export  // switches.export
	);

	wire  [31:0] nios2_data_master_readdata;                           // mm_interconnect_0:NIOS2_data_master_readdata -> NIOS2:d_readdata
	wire         nios2_data_master_waitrequest;                        // mm_interconnect_0:NIOS2_data_master_waitrequest -> NIOS2:d_waitrequest
	wire         nios2_data_master_debugaccess;                        // NIOS2:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:NIOS2_data_master_debugaccess
	wire  [17:0] nios2_data_master_address;                            // NIOS2:d_address -> mm_interconnect_0:NIOS2_data_master_address
	wire   [3:0] nios2_data_master_byteenable;                         // NIOS2:d_byteenable -> mm_interconnect_0:NIOS2_data_master_byteenable
	wire         nios2_data_master_read;                               // NIOS2:d_read -> mm_interconnect_0:NIOS2_data_master_read
	wire         nios2_data_master_write;                              // NIOS2:d_write -> mm_interconnect_0:NIOS2_data_master_write
	wire  [31:0] nios2_data_master_writedata;                          // NIOS2:d_writedata -> mm_interconnect_0:NIOS2_data_master_writedata
	wire  [31:0] nios2_instruction_master_readdata;                    // mm_interconnect_0:NIOS2_instruction_master_readdata -> NIOS2:i_readdata
	wire         nios2_instruction_master_waitrequest;                 // mm_interconnect_0:NIOS2_instruction_master_waitrequest -> NIOS2:i_waitrequest
	wire  [17:0] nios2_instruction_master_address;                     // NIOS2:i_address -> mm_interconnect_0:NIOS2_instruction_master_address
	wire         nios2_instruction_master_read;                        // NIOS2:i_read -> mm_interconnect_0:NIOS2_instruction_master_read
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_chipselect;  // mm_interconnect_0:JTAG_avalon_jtag_slave_chipselect -> JTAG:av_chipselect
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_readdata;    // JTAG:av_readdata -> mm_interconnect_0:JTAG_avalon_jtag_slave_readdata
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest; // JTAG:av_waitrequest -> mm_interconnect_0:JTAG_avalon_jtag_slave_waitrequest
	wire   [0:0] mm_interconnect_0_jtag_avalon_jtag_slave_address;     // mm_interconnect_0:JTAG_avalon_jtag_slave_address -> JTAG:av_address
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_read;        // mm_interconnect_0:JTAG_avalon_jtag_slave_read -> JTAG:av_read_n
	wire         mm_interconnect_0_jtag_avalon_jtag_slave_write;       // mm_interconnect_0:JTAG_avalon_jtag_slave_write -> JTAG:av_write_n
	wire  [31:0] mm_interconnect_0_jtag_avalon_jtag_slave_writedata;   // mm_interconnect_0:JTAG_avalon_jtag_slave_writedata -> JTAG:av_writedata
	wire  [31:0] mm_interconnect_0_sysid_control_slave_readdata;       // SysID:readdata -> mm_interconnect_0:SysID_control_slave_readdata
	wire   [0:0] mm_interconnect_0_sysid_control_slave_address;        // mm_interconnect_0:SysID_control_slave_address -> SysID:address
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_readdata;     // NIOS2:debug_mem_slave_readdata -> mm_interconnect_0:NIOS2_debug_mem_slave_readdata
	wire         mm_interconnect_0_nios2_debug_mem_slave_waitrequest;  // NIOS2:debug_mem_slave_waitrequest -> mm_interconnect_0:NIOS2_debug_mem_slave_waitrequest
	wire         mm_interconnect_0_nios2_debug_mem_slave_debugaccess;  // mm_interconnect_0:NIOS2_debug_mem_slave_debugaccess -> NIOS2:debug_mem_slave_debugaccess
	wire   [8:0] mm_interconnect_0_nios2_debug_mem_slave_address;      // mm_interconnect_0:NIOS2_debug_mem_slave_address -> NIOS2:debug_mem_slave_address
	wire         mm_interconnect_0_nios2_debug_mem_slave_read;         // mm_interconnect_0:NIOS2_debug_mem_slave_read -> NIOS2:debug_mem_slave_read
	wire   [3:0] mm_interconnect_0_nios2_debug_mem_slave_byteenable;   // mm_interconnect_0:NIOS2_debug_mem_slave_byteenable -> NIOS2:debug_mem_slave_byteenable
	wire         mm_interconnect_0_nios2_debug_mem_slave_write;        // mm_interconnect_0:NIOS2_debug_mem_slave_write -> NIOS2:debug_mem_slave_write
	wire  [31:0] mm_interconnect_0_nios2_debug_mem_slave_writedata;    // mm_interconnect_0:NIOS2_debug_mem_slave_writedata -> NIOS2:debug_mem_slave_writedata
	wire         mm_interconnect_0_timercore_s1_chipselect;            // mm_interconnect_0:TimerCore_s1_chipselect -> TimerCore:chipselect
	wire  [15:0] mm_interconnect_0_timercore_s1_readdata;              // TimerCore:readdata -> mm_interconnect_0:TimerCore_s1_readdata
	wire   [2:0] mm_interconnect_0_timercore_s1_address;               // mm_interconnect_0:TimerCore_s1_address -> TimerCore:address
	wire         mm_interconnect_0_timercore_s1_write;                 // mm_interconnect_0:TimerCore_s1_write -> TimerCore:write_n
	wire  [15:0] mm_interconnect_0_timercore_s1_writedata;             // mm_interconnect_0:TimerCore_s1_writedata -> TimerCore:writedata
	wire         mm_interconnect_0_ram_s1_chipselect;                  // mm_interconnect_0:RAM_s1_chipselect -> RAM:chipselect
	wire  [31:0] mm_interconnect_0_ram_s1_readdata;                    // RAM:readdata -> mm_interconnect_0:RAM_s1_readdata
	wire  [12:0] mm_interconnect_0_ram_s1_address;                     // mm_interconnect_0:RAM_s1_address -> RAM:address
	wire   [3:0] mm_interconnect_0_ram_s1_byteenable;                  // mm_interconnect_0:RAM_s1_byteenable -> RAM:byteenable
	wire         mm_interconnect_0_ram_s1_write;                       // mm_interconnect_0:RAM_s1_write -> RAM:write
	wire  [31:0] mm_interconnect_0_ram_s1_writedata;                   // mm_interconnect_0:RAM_s1_writedata -> RAM:writedata
	wire         mm_interconnect_0_ram_s1_clken;                       // mm_interconnect_0:RAM_s1_clken -> RAM:clken
	wire         mm_interconnect_0_segmentsdisplays_s1_chipselect;     // mm_interconnect_0:SegmentsDisplays_s1_chipselect -> SegmentsDisplays:chipselect
	wire  [31:0] mm_interconnect_0_segmentsdisplays_s1_readdata;       // SegmentsDisplays:readdata -> mm_interconnect_0:SegmentsDisplays_s1_readdata
	wire   [1:0] mm_interconnect_0_segmentsdisplays_s1_address;        // mm_interconnect_0:SegmentsDisplays_s1_address -> SegmentsDisplays:address
	wire         mm_interconnect_0_segmentsdisplays_s1_write;          // mm_interconnect_0:SegmentsDisplays_s1_write -> SegmentsDisplays:write_n
	wire  [31:0] mm_interconnect_0_segmentsdisplays_s1_writedata;      // mm_interconnect_0:SegmentsDisplays_s1_writedata -> SegmentsDisplays:writedata
	wire  [31:0] mm_interconnect_0_switches_s1_readdata;               // Switches:readdata -> mm_interconnect_0:Switches_s1_readdata
	wire   [1:0] mm_interconnect_0_switches_s1_address;                // mm_interconnect_0:Switches_s1_address -> Switches:address
	wire  [31:0] mm_interconnect_0_buttons_s1_readdata;                // Buttons:readdata -> mm_interconnect_0:Buttons_s1_readdata
	wire   [1:0] mm_interconnect_0_buttons_s1_address;                 // mm_interconnect_0:Buttons_s1_address -> Buttons:address
	wire         mm_interconnect_0_rom_s1_chipselect;                  // mm_interconnect_0:ROM_s1_chipselect -> ROM:chipselect
	wire  [31:0] mm_interconnect_0_rom_s1_readdata;                    // ROM:readdata -> mm_interconnect_0:ROM_s1_readdata
	wire         mm_interconnect_0_rom_s1_debugaccess;                 // mm_interconnect_0:ROM_s1_debugaccess -> ROM:debugaccess
	wire  [14:0] mm_interconnect_0_rom_s1_address;                     // mm_interconnect_0:ROM_s1_address -> ROM:address
	wire   [3:0] mm_interconnect_0_rom_s1_byteenable;                  // mm_interconnect_0:ROM_s1_byteenable -> ROM:byteenable
	wire         mm_interconnect_0_rom_s1_write;                       // mm_interconnect_0:ROM_s1_write -> ROM:write
	wire  [31:0] mm_interconnect_0_rom_s1_writedata;                   // mm_interconnect_0:ROM_s1_writedata -> ROM:writedata
	wire         mm_interconnect_0_rom_s1_clken;                       // mm_interconnect_0:ROM_s1_clken -> ROM:clken
	wire         mm_interconnect_0_gpioout_s1_chipselect;              // mm_interconnect_0:GpioOut_s1_chipselect -> GpioOut:chipselect
	wire  [31:0] mm_interconnect_0_gpioout_s1_readdata;                // GpioOut:readdata -> mm_interconnect_0:GpioOut_s1_readdata
	wire   [1:0] mm_interconnect_0_gpioout_s1_address;                 // mm_interconnect_0:GpioOut_s1_address -> GpioOut:address
	wire         mm_interconnect_0_gpioout_s1_write;                   // mm_interconnect_0:GpioOut_s1_write -> GpioOut:write_n
	wire  [31:0] mm_interconnect_0_gpioout_s1_writedata;               // mm_interconnect_0:GpioOut_s1_writedata -> GpioOut:writedata
	wire  [31:0] mm_interconnect_0_gpioin_s1_readdata;                 // GpioIn:readdata -> mm_interconnect_0:GpioIn_s1_readdata
	wire   [1:0] mm_interconnect_0_gpioin_s1_address;                  // mm_interconnect_0:GpioIn_s1_address -> GpioIn:address
	wire         mm_interconnect_0_leds_s1_chipselect;                 // mm_interconnect_0:Leds_s1_chipselect -> Leds:chipselect
	wire  [31:0] mm_interconnect_0_leds_s1_readdata;                   // Leds:readdata -> mm_interconnect_0:Leds_s1_readdata
	wire   [1:0] mm_interconnect_0_leds_s1_address;                    // mm_interconnect_0:Leds_s1_address -> Leds:address
	wire         mm_interconnect_0_leds_s1_write;                      // mm_interconnect_0:Leds_s1_write -> Leds:write_n
	wire  [31:0] mm_interconnect_0_leds_s1_writedata;                  // mm_interconnect_0:Leds_s1_writedata -> Leds:writedata
	wire         irq_mapper_receiver0_irq;                             // TimerCore:irq -> irq_mapper:receiver0_irq
	wire         irq_mapper_receiver1_irq;                             // JTAG:av_irq -> irq_mapper:receiver1_irq
	wire  [31:0] nios2_irq_irq;                                        // irq_mapper:sender_irq -> NIOS2:irq
	wire         rst_controller_reset_out_reset;                       // rst_controller:reset_out -> [Buttons:reset_n, GpioIn:reset_n, GpioOut:reset_n, JTAG:rst_n, Leds:reset_n, NIOS2:reset_n, RAM:reset, ROM:reset, SegmentsDisplays:reset_n, Switches:reset_n, SysID:reset_n, TimerCore:reset_n, irq_mapper:reset, mm_interconnect_0:NIOS2_reset_reset_bridge_in_reset_reset, rst_translator:in_reset]
	wire         rst_controller_reset_out_reset_req;                   // rst_controller:reset_req -> [NIOS2:reset_req, RAM:reset_req, ROM:reset_req, rst_translator:reset_req_in]
	wire         nios2_debug_reset_request_reset;                      // NIOS2:debug_reset_request -> rst_controller:reset_in1

	TimerSoC_Buttons buttons (
		.clk      (clk_clk),                               //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),       //               reset.reset_n
		.address  (mm_interconnect_0_buttons_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_buttons_s1_readdata), //                    .readdata
		.in_port  (buttons_export)                         // external_connection.export
	);

	TimerSoC_GpioIn gpioin (
		.clk      (clk_clk),                              //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address  (mm_interconnect_0_gpioin_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_gpioin_s1_readdata), //                    .readdata
		.in_port  (gpio_in_export)                        // external_connection.export
	);

	TimerSoC_GpioOut gpioout (
		.clk        (clk_clk),                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),         //               reset.reset_n
		.address    (mm_interconnect_0_gpioout_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_gpioout_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_gpioout_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_gpioout_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_gpioout_s1_readdata),   //                    .readdata
		.out_port   (gpio_out_export)                          // external_connection.export
	);

	TimerSoC_JTAG jtag (
		.clk            (clk_clk),                                              //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                      //             reset.reset_n
		.av_chipselect  (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //                  .address
		.av_read_n      (~mm_interconnect_0_jtag_avalon_jtag_slave_read),       //                  .read_n
		.av_readdata    (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                  .readdata
		.av_write_n     (~mm_interconnect_0_jtag_avalon_jtag_slave_write),      //                  .write_n
		.av_writedata   (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                  .writedata
		.av_waitrequest (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver1_irq)                              //               irq.irq
	);

	TimerSoC_Leds leds (
		.clk        (clk_clk),                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),      //               reset.reset_n
		.address    (mm_interconnect_0_leds_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_leds_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_leds_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_leds_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_leds_s1_readdata),   //                    .readdata
		.out_port   (leds_export)                           // external_connection.export
	);

	TimerSoC_NIOS2 nios2 (
		.clk                                 (clk_clk),                                             //                       clk.clk
		.reset_n                             (~rst_controller_reset_out_reset),                     //                     reset.reset_n
		.reset_req                           (rst_controller_reset_out_reset_req),                  //                          .reset_req
		.d_address                           (nios2_data_master_address),                           //               data_master.address
		.d_byteenable                        (nios2_data_master_byteenable),                        //                          .byteenable
		.d_read                              (nios2_data_master_read),                              //                          .read
		.d_readdata                          (nios2_data_master_readdata),                          //                          .readdata
		.d_waitrequest                       (nios2_data_master_waitrequest),                       //                          .waitrequest
		.d_write                             (nios2_data_master_write),                             //                          .write
		.d_writedata                         (nios2_data_master_writedata),                         //                          .writedata
		.debug_mem_slave_debugaccess_to_roms (nios2_data_master_debugaccess),                       //                          .debugaccess
		.i_address                           (nios2_instruction_master_address),                    //        instruction_master.address
		.i_read                              (nios2_instruction_master_read),                       //                          .read
		.i_readdata                          (nios2_instruction_master_readdata),                   //                          .readdata
		.i_waitrequest                       (nios2_instruction_master_waitrequest),                //                          .waitrequest
		.irq                                 (nios2_irq_irq),                                       //                       irq.irq
		.debug_reset_request                 (nios2_debug_reset_request_reset),                     //       debug_reset_request.reset
		.debug_mem_slave_address             (mm_interconnect_0_nios2_debug_mem_slave_address),     //           debug_mem_slave.address
		.debug_mem_slave_byteenable          (mm_interconnect_0_nios2_debug_mem_slave_byteenable),  //                          .byteenable
		.debug_mem_slave_debugaccess         (mm_interconnect_0_nios2_debug_mem_slave_debugaccess), //                          .debugaccess
		.debug_mem_slave_read                (mm_interconnect_0_nios2_debug_mem_slave_read),        //                          .read
		.debug_mem_slave_readdata            (mm_interconnect_0_nios2_debug_mem_slave_readdata),    //                          .readdata
		.debug_mem_slave_waitrequest         (mm_interconnect_0_nios2_debug_mem_slave_waitrequest), //                          .waitrequest
		.debug_mem_slave_write               (mm_interconnect_0_nios2_debug_mem_slave_write),       //                          .write
		.debug_mem_slave_writedata           (mm_interconnect_0_nios2_debug_mem_slave_writedata),   //                          .writedata
		.dummy_ci_port                       ()                                                     // custom_instruction_master.readra
	);

	TimerSoC_RAM ram (
		.clk        (clk_clk),                             //   clk1.clk
		.address    (mm_interconnect_0_ram_s1_address),    //     s1.address
		.clken      (mm_interconnect_0_ram_s1_clken),      //       .clken
		.chipselect (mm_interconnect_0_ram_s1_chipselect), //       .chipselect
		.write      (mm_interconnect_0_ram_s1_write),      //       .write
		.readdata   (mm_interconnect_0_ram_s1_readdata),   //       .readdata
		.writedata  (mm_interconnect_0_ram_s1_writedata),  //       .writedata
		.byteenable (mm_interconnect_0_ram_s1_byteenable), //       .byteenable
		.reset      (rst_controller_reset_out_reset),      // reset1.reset
		.reset_req  (rst_controller_reset_out_reset_req),  //       .reset_req
		.freeze     (1'b0)                                 // (terminated)
	);

	TimerSoC_ROM rom (
		.clk         (clk_clk),                              //   clk1.clk
		.address     (mm_interconnect_0_rom_s1_address),     //     s1.address
		.debugaccess (mm_interconnect_0_rom_s1_debugaccess), //       .debugaccess
		.clken       (mm_interconnect_0_rom_s1_clken),       //       .clken
		.chipselect  (mm_interconnect_0_rom_s1_chipselect),  //       .chipselect
		.write       (mm_interconnect_0_rom_s1_write),       //       .write
		.readdata    (mm_interconnect_0_rom_s1_readdata),    //       .readdata
		.writedata   (mm_interconnect_0_rom_s1_writedata),   //       .writedata
		.byteenable  (mm_interconnect_0_rom_s1_byteenable),  //       .byteenable
		.reset       (rst_controller_reset_out_reset),       // reset1.reset
		.reset_req   (rst_controller_reset_out_reset_req),   //       .reset_req
		.freeze      (1'b0)                                  // (terminated)
	);

	TimerSoC_SegmentsDisplays segmentsdisplays (
		.clk        (clk_clk),                                          //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                  //               reset.reset_n
		.address    (mm_interconnect_0_segmentsdisplays_s1_address),    //                  s1.address
		.write_n    (~mm_interconnect_0_segmentsdisplays_s1_write),     //                    .write_n
		.writedata  (mm_interconnect_0_segmentsdisplays_s1_writedata),  //                    .writedata
		.chipselect (mm_interconnect_0_segmentsdisplays_s1_chipselect), //                    .chipselect
		.readdata   (mm_interconnect_0_segmentsdisplays_s1_readdata),   //                    .readdata
		.out_port   (displays_export)                                   // external_connection.export
	);

	TimerSoC_Buttons switches (
		.clk      (clk_clk),                                //                 clk.clk
		.reset_n  (~rst_controller_reset_out_reset),        //               reset.reset_n
		.address  (mm_interconnect_0_switches_s1_address),  //                  s1.address
		.readdata (mm_interconnect_0_switches_s1_readdata), //                    .readdata
		.in_port  (switches_export)                         // external_connection.export
	);

	TimerSoC_SysID sysid (
		.clock    (clk_clk),                                        //           clk.clk
		.reset_n  (~rst_controller_reset_out_reset),                //         reset.reset_n
		.readdata (mm_interconnect_0_sysid_control_slave_readdata), // control_slave.readdata
		.address  (mm_interconnect_0_sysid_control_slave_address)   //              .address
	);

	TimerSoC_TimerCore timercore (
		.clk        (clk_clk),                                   //   clk.clk
		.reset_n    (~rst_controller_reset_out_reset),           // reset.reset_n
		.address    (mm_interconnect_0_timercore_s1_address),    //    s1.address
		.writedata  (mm_interconnect_0_timercore_s1_writedata),  //      .writedata
		.readdata   (mm_interconnect_0_timercore_s1_readdata),   //      .readdata
		.chipselect (mm_interconnect_0_timercore_s1_chipselect), //      .chipselect
		.write_n    (~mm_interconnect_0_timercore_s1_write),     //      .write_n
		.irq        (irq_mapper_receiver0_irq)                   //   irq.irq
	);

	TimerSoC_mm_interconnect_0 mm_interconnect_0 (
		.Clock_clk_clk                           (clk_clk),                                              //                         Clock_clk.clk
		.NIOS2_reset_reset_bridge_in_reset_reset (rst_controller_reset_out_reset),                       // NIOS2_reset_reset_bridge_in_reset.reset
		.NIOS2_data_master_address               (nios2_data_master_address),                            //                 NIOS2_data_master.address
		.NIOS2_data_master_waitrequest           (nios2_data_master_waitrequest),                        //                                  .waitrequest
		.NIOS2_data_master_byteenable            (nios2_data_master_byteenable),                         //                                  .byteenable
		.NIOS2_data_master_read                  (nios2_data_master_read),                               //                                  .read
		.NIOS2_data_master_readdata              (nios2_data_master_readdata),                           //                                  .readdata
		.NIOS2_data_master_write                 (nios2_data_master_write),                              //                                  .write
		.NIOS2_data_master_writedata             (nios2_data_master_writedata),                          //                                  .writedata
		.NIOS2_data_master_debugaccess           (nios2_data_master_debugaccess),                        //                                  .debugaccess
		.NIOS2_instruction_master_address        (nios2_instruction_master_address),                     //          NIOS2_instruction_master.address
		.NIOS2_instruction_master_waitrequest    (nios2_instruction_master_waitrequest),                 //                                  .waitrequest
		.NIOS2_instruction_master_read           (nios2_instruction_master_read),                        //                                  .read
		.NIOS2_instruction_master_readdata       (nios2_instruction_master_readdata),                    //                                  .readdata
		.Buttons_s1_address                      (mm_interconnect_0_buttons_s1_address),                 //                        Buttons_s1.address
		.Buttons_s1_readdata                     (mm_interconnect_0_buttons_s1_readdata),                //                                  .readdata
		.GpioIn_s1_address                       (mm_interconnect_0_gpioin_s1_address),                  //                         GpioIn_s1.address
		.GpioIn_s1_readdata                      (mm_interconnect_0_gpioin_s1_readdata),                 //                                  .readdata
		.GpioOut_s1_address                      (mm_interconnect_0_gpioout_s1_address),                 //                        GpioOut_s1.address
		.GpioOut_s1_write                        (mm_interconnect_0_gpioout_s1_write),                   //                                  .write
		.GpioOut_s1_readdata                     (mm_interconnect_0_gpioout_s1_readdata),                //                                  .readdata
		.GpioOut_s1_writedata                    (mm_interconnect_0_gpioout_s1_writedata),               //                                  .writedata
		.GpioOut_s1_chipselect                   (mm_interconnect_0_gpioout_s1_chipselect),              //                                  .chipselect
		.JTAG_avalon_jtag_slave_address          (mm_interconnect_0_jtag_avalon_jtag_slave_address),     //            JTAG_avalon_jtag_slave.address
		.JTAG_avalon_jtag_slave_write            (mm_interconnect_0_jtag_avalon_jtag_slave_write),       //                                  .write
		.JTAG_avalon_jtag_slave_read             (mm_interconnect_0_jtag_avalon_jtag_slave_read),        //                                  .read
		.JTAG_avalon_jtag_slave_readdata         (mm_interconnect_0_jtag_avalon_jtag_slave_readdata),    //                                  .readdata
		.JTAG_avalon_jtag_slave_writedata        (mm_interconnect_0_jtag_avalon_jtag_slave_writedata),   //                                  .writedata
		.JTAG_avalon_jtag_slave_waitrequest      (mm_interconnect_0_jtag_avalon_jtag_slave_waitrequest), //                                  .waitrequest
		.JTAG_avalon_jtag_slave_chipselect       (mm_interconnect_0_jtag_avalon_jtag_slave_chipselect),  //                                  .chipselect
		.Leds_s1_address                         (mm_interconnect_0_leds_s1_address),                    //                           Leds_s1.address
		.Leds_s1_write                           (mm_interconnect_0_leds_s1_write),                      //                                  .write
		.Leds_s1_readdata                        (mm_interconnect_0_leds_s1_readdata),                   //                                  .readdata
		.Leds_s1_writedata                       (mm_interconnect_0_leds_s1_writedata),                  //                                  .writedata
		.Leds_s1_chipselect                      (mm_interconnect_0_leds_s1_chipselect),                 //                                  .chipselect
		.NIOS2_debug_mem_slave_address           (mm_interconnect_0_nios2_debug_mem_slave_address),      //             NIOS2_debug_mem_slave.address
		.NIOS2_debug_mem_slave_write             (mm_interconnect_0_nios2_debug_mem_slave_write),        //                                  .write
		.NIOS2_debug_mem_slave_read              (mm_interconnect_0_nios2_debug_mem_slave_read),         //                                  .read
		.NIOS2_debug_mem_slave_readdata          (mm_interconnect_0_nios2_debug_mem_slave_readdata),     //                                  .readdata
		.NIOS2_debug_mem_slave_writedata         (mm_interconnect_0_nios2_debug_mem_slave_writedata),    //                                  .writedata
		.NIOS2_debug_mem_slave_byteenable        (mm_interconnect_0_nios2_debug_mem_slave_byteenable),   //                                  .byteenable
		.NIOS2_debug_mem_slave_waitrequest       (mm_interconnect_0_nios2_debug_mem_slave_waitrequest),  //                                  .waitrequest
		.NIOS2_debug_mem_slave_debugaccess       (mm_interconnect_0_nios2_debug_mem_slave_debugaccess),  //                                  .debugaccess
		.RAM_s1_address                          (mm_interconnect_0_ram_s1_address),                     //                            RAM_s1.address
		.RAM_s1_write                            (mm_interconnect_0_ram_s1_write),                       //                                  .write
		.RAM_s1_readdata                         (mm_interconnect_0_ram_s1_readdata),                    //                                  .readdata
		.RAM_s1_writedata                        (mm_interconnect_0_ram_s1_writedata),                   //                                  .writedata
		.RAM_s1_byteenable                       (mm_interconnect_0_ram_s1_byteenable),                  //                                  .byteenable
		.RAM_s1_chipselect                       (mm_interconnect_0_ram_s1_chipselect),                  //                                  .chipselect
		.RAM_s1_clken                            (mm_interconnect_0_ram_s1_clken),                       //                                  .clken
		.ROM_s1_address                          (mm_interconnect_0_rom_s1_address),                     //                            ROM_s1.address
		.ROM_s1_write                            (mm_interconnect_0_rom_s1_write),                       //                                  .write
		.ROM_s1_readdata                         (mm_interconnect_0_rom_s1_readdata),                    //                                  .readdata
		.ROM_s1_writedata                        (mm_interconnect_0_rom_s1_writedata),                   //                                  .writedata
		.ROM_s1_byteenable                       (mm_interconnect_0_rom_s1_byteenable),                  //                                  .byteenable
		.ROM_s1_chipselect                       (mm_interconnect_0_rom_s1_chipselect),                  //                                  .chipselect
		.ROM_s1_clken                            (mm_interconnect_0_rom_s1_clken),                       //                                  .clken
		.ROM_s1_debugaccess                      (mm_interconnect_0_rom_s1_debugaccess),                 //                                  .debugaccess
		.SegmentsDisplays_s1_address             (mm_interconnect_0_segmentsdisplays_s1_address),        //               SegmentsDisplays_s1.address
		.SegmentsDisplays_s1_write               (mm_interconnect_0_segmentsdisplays_s1_write),          //                                  .write
		.SegmentsDisplays_s1_readdata            (mm_interconnect_0_segmentsdisplays_s1_readdata),       //                                  .readdata
		.SegmentsDisplays_s1_writedata           (mm_interconnect_0_segmentsdisplays_s1_writedata),      //                                  .writedata
		.SegmentsDisplays_s1_chipselect          (mm_interconnect_0_segmentsdisplays_s1_chipselect),     //                                  .chipselect
		.Switches_s1_address                     (mm_interconnect_0_switches_s1_address),                //                       Switches_s1.address
		.Switches_s1_readdata                    (mm_interconnect_0_switches_s1_readdata),               //                                  .readdata
		.SysID_control_slave_address             (mm_interconnect_0_sysid_control_slave_address),        //               SysID_control_slave.address
		.SysID_control_slave_readdata            (mm_interconnect_0_sysid_control_slave_readdata),       //                                  .readdata
		.TimerCore_s1_address                    (mm_interconnect_0_timercore_s1_address),               //                      TimerCore_s1.address
		.TimerCore_s1_write                      (mm_interconnect_0_timercore_s1_write),                 //                                  .write
		.TimerCore_s1_readdata                   (mm_interconnect_0_timercore_s1_readdata),              //                                  .readdata
		.TimerCore_s1_writedata                  (mm_interconnect_0_timercore_s1_writedata),             //                                  .writedata
		.TimerCore_s1_chipselect                 (mm_interconnect_0_timercore_s1_chipselect)             //                                  .chipselect
	);

	TimerSoC_irq_mapper irq_mapper (
		.clk           (clk_clk),                        //       clk.clk
		.reset         (rst_controller_reset_out_reset), // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq),       // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq),       // receiver1.irq
		.sender_irq    (nios2_irq_irq)                   //    sender.irq
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS          (2),
		.OUTPUT_RESET_SYNC_EDGES   ("deassert"),
		.SYNC_DEPTH                (2),
		.RESET_REQUEST_PRESENT     (1),
		.RESET_REQ_WAIT_TIME       (1),
		.MIN_RST_ASSERTION_TIME    (3),
		.RESET_REQ_EARLY_DSRT_TIME (1),
		.USE_RESET_REQUEST_IN0     (0),
		.USE_RESET_REQUEST_IN1     (0),
		.USE_RESET_REQUEST_IN2     (0),
		.USE_RESET_REQUEST_IN3     (0),
		.USE_RESET_REQUEST_IN4     (0),
		.USE_RESET_REQUEST_IN5     (0),
		.USE_RESET_REQUEST_IN6     (0),
		.USE_RESET_REQUEST_IN7     (0),
		.USE_RESET_REQUEST_IN8     (0),
		.USE_RESET_REQUEST_IN9     (0),
		.USE_RESET_REQUEST_IN10    (0),
		.USE_RESET_REQUEST_IN11    (0),
		.USE_RESET_REQUEST_IN12    (0),
		.USE_RESET_REQUEST_IN13    (0),
		.USE_RESET_REQUEST_IN14    (0),
		.USE_RESET_REQUEST_IN15    (0),
		.ADAPT_RESET_REQUEST       (0)
	) rst_controller (
		.reset_in0      (~reset_reset_n),                     // reset_in0.reset
		.reset_in1      (nios2_debug_reset_request_reset),    // reset_in1.reset
		.clk            (clk_clk),                            //       clk.clk
		.reset_out      (rst_controller_reset_out_reset),     // reset_out.reset
		.reset_req      (rst_controller_reset_out_reset_req), //          .reset_req
		.reset_req_in0  (1'b0),                               // (terminated)
		.reset_req_in1  (1'b0),                               // (terminated)
		.reset_in2      (1'b0),                               // (terminated)
		.reset_req_in2  (1'b0),                               // (terminated)
		.reset_in3      (1'b0),                               // (terminated)
		.reset_req_in3  (1'b0),                               // (terminated)
		.reset_in4      (1'b0),                               // (terminated)
		.reset_req_in4  (1'b0),                               // (terminated)
		.reset_in5      (1'b0),                               // (terminated)
		.reset_req_in5  (1'b0),                               // (terminated)
		.reset_in6      (1'b0),                               // (terminated)
		.reset_req_in6  (1'b0),                               // (terminated)
		.reset_in7      (1'b0),                               // (terminated)
		.reset_req_in7  (1'b0),                               // (terminated)
		.reset_in8      (1'b0),                               // (terminated)
		.reset_req_in8  (1'b0),                               // (terminated)
		.reset_in9      (1'b0),                               // (terminated)
		.reset_req_in9  (1'b0),                               // (terminated)
		.reset_in10     (1'b0),                               // (terminated)
		.reset_req_in10 (1'b0),                               // (terminated)
		.reset_in11     (1'b0),                               // (terminated)
		.reset_req_in11 (1'b0),                               // (terminated)
		.reset_in12     (1'b0),                               // (terminated)
		.reset_req_in12 (1'b0),                               // (terminated)
		.reset_in13     (1'b0),                               // (terminated)
		.reset_req_in13 (1'b0),                               // (terminated)
		.reset_in14     (1'b0),                               // (terminated)
		.reset_req_in14 (1'b0),                               // (terminated)
		.reset_in15     (1'b0),                               // (terminated)
		.reset_req_in15 (1'b0)                                // (terminated)
	);

endmodule
